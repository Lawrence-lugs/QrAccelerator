// ROM for microcode looper

import qracc_pkg::*;

module ucode_ctrl #(
    parameter dataWidth = 32,
    parameter addrWidth = 32
) (
    input [dataWidth-1:0] addr,
    output [dataWidth-1:0] idx
);



endmodule