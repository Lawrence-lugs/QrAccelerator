`ifndef PARAMETERS_FILE
`define PARAMETERS_FILE
`define PYTEST_GENERATED_PARAMS
`define PYTEST_GENERATED_PARAMS
`define SRAM_ROWS 256
`define SRAM_COLS 256
`define QRACC_INPUT_BITS 8
`define QRACC_OUTPUT_BITS 8
`define GB_INT_IF_WIDTH 256
`define NODUMP 1
`define NOTPLITZTRACK 1
`define NOIOFILES 1
`define SNOOP_OFMAP 1
`define TRACK_STATISTICS 1
`endif // PARAMETERS_FILE
