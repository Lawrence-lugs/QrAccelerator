// Overall controller for QRAcc
// Microcode looper

module qracc_control #(

) (
    input clk, nrst,
    input qracc_start_i,
    input loop_config_t loop_config

    // Outputs
);

// Parameters


// Signals
logic [31:0] pc;
logic jump;
logic [31:0] jump_addr;

// Modules




endmodule