`ifndef PARAMETERS_FILE
`define PARAMETERS_FILE
`define PYTEST_GENERATED_PARAMS
`define PYTEST_GENERATED_PARAMS
`define SRAM_ROWS 256
`define SRAM_COLS 256
`define QRACC_INPUT_BITS 8
`define QRACC_OUTPUT_BITS 8
`define GB_INT_IF_WIDTH 256
`define FILTER_SIZE_X 3
`define FILTER_SIZE_Y 3
`define OFMAP_SIZE 65536
`define IFMAP_SIZE 8748
`define IFMAP_DIMX 16
`define IFMAP_DIMY 16
`define OFMAP_DIMX 16
`define OFMAP_DIMY 16
`define IN_CHANNELS 27
`define OUT_CHANNELS 256
`define MAPPED_MATRIX_OFFSET_X 0
`define MAPPED_MATRIX_OFFSET_Y 0
`define STRIDE_X 1
`define STRIDE_Y 1
`define UNSIGNED_ACTS 1
`define NUM_ADC_REF_RANGE_SHIFTS 4
`endif // PARAMETERS_FILE
