qracc_pkg.svh