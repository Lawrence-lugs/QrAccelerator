`timescale 1ns/1ps

package qracc_pkg;

    parameter numRows = 128;
    parameter numCols = 32;
    parameter numAdcBits = 4;
    parameter compCount = (2**numAdcBits)-1;
    parameter numCfgBits = 8;

    typedef struct packed {        
        logic [numCfgBits-1:0] n_input_bits_cfg;
        // logic [numCfgBits-1:0] n_adc_bits_cfg;
        logic binary_cfg;
    } qracc_config_t;

    typedef struct {
        // SWITCH MATRIX
        logic [numRows-1:0] VDR_SEL;
        logic [numRows-1:0] VDR_SELB;
        logic [numRows-1:0] VSS_SEL;
        logic [numRows-1:0] VSS_SELB;
        logic [numRows-1:0] VRST_SEL;
        logic [numRows-1:0] VRST_SELB;

        // SRAM
        logic [numRows-1:0] WL;
        logic PCH;
        logic [numCols-1:0] WR_DATA;
        logic WRITE;
        logic [numCols-1:0] CSEL;
        logic SAEN;

        // ADC
        logic NF;
        logic NFB;
        logic M2A;
        logic M2AB;
        logic R2A;
        logic R2AB;

        // Clock
        logic CLK;
    } to_analog_t;

    typedef struct {
        logic [numCols-1:0] SA_OUT;
        logic [compCount*numCols-1:0] ADC_OUT;
    } from_analog_t;

endpackage