`ifndef PARAMETERS_FILE
`define PARAMETERS_FILE
`define PYTEST_GENERATED_PARAMS
`define PYTEST_GENERATED_PARAMS
`define SRAM_ROWS 256
`define SRAM_COLS 32
`define QRACC_INPUT_BITS 8
`define QRACC_OUTPUT_BITS 8
`define GB_INT_IF_WIDTH 2048
`define FILTER_SIZE_X 3
`define FILTER_SIZE_Y 3
`define OFMAP_SIZE 32768
`define IFMAP_SIZE 3468
`define IFMAP_DIMX 34
`define IFMAP_DIMY 34
`define OFMAP_DIMX 32
`define OFMAP_DIMY 32
`define IN_CHANNELS 3
`define OUT_CHANNELS 32
`define MAPPED_MATRIX_OFFSET_X 0
`define MAPPED_MATRIX_OFFSET_Y 0
`define UNSIGNED_ACTS 1
`endif // PARAMETERS_FILE
