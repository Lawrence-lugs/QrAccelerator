../../../c3sram_periphery/rtl/c3sram_mac_wrap.sv