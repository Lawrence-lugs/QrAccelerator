/home/lquizon/lawrence-workspace/sram_interface/rtl/sram_32bank_8b.sv