`define SRAM_ROWS 256
`define SRAM_COLS 32
`define QRACC_INPUT_BITS 8
`define QRACC_OUTPUT_BITS 8
`define GB_INT_IF_WIDTH 2048
`define FILTER_SIZE_X 3
`define FILTER_SIZE_Y 3
`define OFMAP_SIZE 16
`define IFMAP_SIZE 972
`define IFMAP_DIMX 18
`define IFMAP_DIMY 18
`define OFMAP_DIMX 16
`define OFMAP_DIMY 16
`define IN_CHANNELS 3
`define OUT_CHANNELS 32
`define MAPPED_MATRIX_OFFSET_X 0
`define MAPPED_MATRIX_OFFSET_Y 0
