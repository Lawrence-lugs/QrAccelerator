`define SRAM_ROWS 256
`define SRAM_COLS 32
`define QRACC_INPUT_BITS 4
`define QRACC_OUTPUT_BITS 4
`define GB_INT_IF_WIDTH 1024
